module imem (
	input  [ 7:0] addr,
	output [31:0] data
);

	reg [31:0] data;

	// r6 ith element
	// r1 index
	// r2 sum
	// r3 n (gp)
	// r5 address of ith element
	// r10 address of sum (gp +4)

	always @(addr) begin
		case(addr)
			//  addi r1 r0 0
			// op- 001000
			// rs- 00000
			// rt- 00001
			// i- 0000 0000 0000 0000
			00 : data = 32'b00100000000000010000000000000000;

			// addi r2 r0 0
			// op- 001000
			// rs- 00000
			// rt- 00010
			// i- 0000 0000 0000 0000
			04 : data = 32'b00100000000000100000000000000000;

			// addi r4 $gp 0
			// op- 001000
			// rt- 00100
			// rs- 11000
			// i-  0000 0000 0000 0000
			08 : data = 32'b00100011000001000000000000000000;

			// lw r3 r4
			// op- 100011
			// rt- 00011
			// rs- 00100
			// i- 0000 0000 0000 0000
			12 : data = 32'b10001100100000110000000000000000;

			// addi r5 $gp 8
			// op- 001000
			// rt- 00101
			// rs- 11000
			// i- 0000 0000 0000 1000
			16 : data = 32'b00100011000001010000000000001000;

			// addi r10 $gp 4
			// op- 001000
			// rt- 01010
			// rs- 11000
			// i-  0000 0000 0000 0100
			20 : data = 32'b00100011000010100000000000000100;

			// beq r1 r3 end
			// op- 000100
			// rs - 00001
			// rt - 00011
			// im - end-here-4
			24 : data = 32'b00010000001000110000000000000101;

			// lw r6 r5 0 
			// op-100011
			// rs-00101
			// rt-00110
			// i - 0
			28 : data = 32'b10001100101001100000000000000000;

			// add r2 r2 r6
			// op- 000000
			// rd- - 00010
			// rs - 00010
			// rt - 00110
			// shamt  - 00000
			// funct - 100000
			32 : data = 32'b00000000010001100001000000100000;

			// addi r5 r5 4
			// op - 001000
			// rt - 000101
			// rs - 000101
			// im - 4
			36 : data = 32'b00100000101001010000000000000100;

			//addi r1 r1 1
			// op - 001000
			// rt - 00001
			// rs - 00001
			// im - 00000000000000001
			40 : data = 32'b00100000001000010000000000000001;

			// j start 
			// op - 000010
			// addr - start
			// 000010 000000000000000000110
			44 : data = 32'b00001000000000000000000000000110;

			//sw r10 r6
			// op - 101011
			// rs - 01010
			// rt - 00010
			// imm - 0
			48 : data = 32'b10101101010000100000000000000000;

			// addi r4 r0 10 (argument for syscall)
			// op- 001000
			// rs- 00000
			// rt- 00100
			// i- 0000 0000 0000 1010
			52 : data = 32'b00100000000001000000000000001010;

			// syscall
			// op - 001100
			56 : data = 32'b00110000000000000000000000000000;
		endcase
	end
endmodule
